library ieee;
use ieee.numeric_std.all;

package common is
  subtype word is unsigned(7 downto 0);
end package common;

