library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.std_logic_unsigned.all;
use ieee.numeric_std.all;
library lcd;
use lcd.LCDCommunication.all;
use lcd.LCDInterrupt.all;

entity LCD_Controller is
    Port ( 
		iclock 		  : in std_logic;
		userControl   : in UserControl;
		lcdInterrupt  : out LCdInterrupt;--H: busy L: Ready
		lcdControl    : out LCDControl);
end LCD_Controller;

architecture Behavioral of LCD_Controller is

component Wait_Timer is
    Generic( 
           Board_Clock : INTEGER := 125_000_000);--ns
    Port ( 
           iclk : in STD_LOGIC;
           ienable : in STD_LOGIC;
           iwait_time : in INTEGER;--in ns
           oenable : out STD_LOGIC);
end component;
		
	type ModeStates is (Power_Up_Mode, Initialize_Mode, User_Mode); --All Modes

	constant power_up_time				: integer := 20_000_000;--20 ms
	constant enable_time           		: integer := 5_000_000;--5ms (15 ms period for enable pulse)
	constant initialize_instructions    : integer := 13;--que

	signal internal_enable_state		: integer range 0 to 2;
	signal time_counter					: integer := 0;
	signal Mode 						: ModeStates := Power_Up_Mode;
	signal initialize_state			    : integer range 0 to initialize_instructions;--one extra int value for change
	signal Data_s						: unsigned(7 downto 0);
    --wait timmer signals
    signal oenable_s : STD_LOGIC := '0';
    signal ienable_s : STD_LOGIC := '0';
    signal iwait_time_s : INTEGER := 0;--in ns
    
begin
    
    enable_pulse : process(iclock)--and wait time for power up
    begin
    case Mode is
        when Power_Up_Mode =>
            iwait_time_s <= power_up_time;--20ms
            ienable_s <= '1';
            if oenable_s = '1' then
                ienable_s <= '0';
            end if;
        when Initialize_Mode =>
             iwait_time_s <= enable_time;--5ms
             ienable_s <= '1';
             if oenable_s = '1' then
                 ienable_s <= '0';
             end if;
        when others =>
    end case;
    end process;
    
    Mode_Changes : process(iclock)
    begin
    case Mode is
        when Power_Up_Mode =>
            if oenable_s = '1' then
                Mode <= Initialize_Mode;
            end if;
        when Initialize_Mode =>
            if initialize_state = initialize_instructions AND internal_enable_state = 0 then
                Mode <= User_Mode;
            end if;
        when User_Mode =>
            if userControl.Reset = '1' then
                Mode <= Initialize_Mode;
            end if;
    end case;
    end process;
    
    with initialize_state select
        Data_s <=
            X"3" when 0,--8 bit interface
            X"3" when 1,
            X"3" when 2,
            X"2" when 3,--4 bit interface
            "0010" when 4,
            "1XXX" when 5,-- function set number of lines: 2
            "0000" when 6,
            "1000" when 7,--Display, cursor, Blinking off
            "0000" when 8,
            "0001" when 9,--clear display
            "0000" when 10,
            "0110" when 11,--inc cursor to the right when writing and dont shift screen
            "0000" when 12,
            "1100" when 13;--Display on
        
    process(iclock, Mode, internal_enable_state)--Mode process
    begin
    if rising_edge(iclock) then
        case Mode is
            when Power_Up_Mode =>
                lcdControl.RS			<= '0';
                lcdControl.RW			<= '0';
                lcdInterrupt.isBusy		<= '1';
                lcdControl.enable 	    <= '0';
                lcdControl.nibble 		<= X"28";
            when Initialize_Mode =>
                lcdControl.nibble 		<= Data_s;
                lcdControl.RS			<= '0';
                lcdControl.RW			<= '0';
                lcdInterrupt.isBusy		<= '1';
                case internal_enable_state is
                    when 0 => 	
                        lcdControl.enable <= '0';
                    when 1 =>
                        lcdControl.enable <= '1';
                    when 2 =>
                        lcdControl.enable <= '0';			
                end case;
                if oenable_s = '1' then
                    if internal_enable_state < 2 then
                         internal_enable_state <= internal_enable_state + 1;
                     else
                         internal_enable_state <= 0;
                     end if;
                end if; 
            when User_Mode =>
                lcdControl.nibble 		<= UserControl.nibble;
                lcdControl.RS			<= UserControl.RS;
                lcdControl.RW			<= '0';
                lcdInterrupt.isBusy		<= '0';
                lcdControl.enable 	    <= UserControl.enable;
        end case;
    end if;
    end process;

Inst_Wait_Timer : Wait_Timer
    Generic Map ( 
           Board_Clock => 125_000_000)--ns
    Port Map ( 
           iclk => iclock,
           ienable => ienable_s,
           iwait_time => iwait_time_s,
           oenable => oenable_s);
end Behavioral;